// flappy_bird_control.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module flappy_bird_control (
		output wire [15:0] bird_x_export_export,             //             bird_x_export.export
		output wire [15:0] bird_y2_export_export,            //            bird_y2_export.export
		output wire [15:0] bird_y_export_export,             //             bird_y_export.export
		input  wire        clk_clk,                          //                       clk.clk
		output wire [15:0] first2_export_export,             //             first2_export.export
		output wire [15:0] first_export_export,              //              first_export.export
		input  wire [7:0]  keycode_export_export,            //            keycode_export.export
		output wire [15:0] level_external_connection_export, // level_external_connection.export
		output wire [15:0] pipe1_export_export,              //              pipe1_export.export
		output wire [15:0] pipe2_export_export,              //              pipe2_export.export
		output wire [15:0] pipe3_export_export,              //              pipe3_export.export
		output wire [15:0] pipe4_export_export,              //              pipe4_export.export
		output wire [15:0] pipe5_export_export,              //              pipe5_export.export
		output wire [15:0] pipe_x_export_export,             //             pipe_x_export.export
		input  wire        press_export_export,              //              press_export.export
		input  wire        reset_reset_n,                    //                     reset.reset_n
		output wire [15:0] scorex2_export_export,            //            scorex2_export.export
		output wire [15:0] scorex_export_export,             //             scorex_export.export
		output wire [15:0] scorey2_export_export,            //            scorey2_export.export
		output wire [15:0] scorey_export_export,             //             scorey_export.export
		output wire        sdram_clk_clk,                    //                 sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                  //                sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                    //                          .ba
		output wire        sdram_wire_cas_n,                 //                          .cas_n
		output wire        sdram_wire_cke,                   //                          .cke
		output wire        sdram_wire_cs_n,                  //                          .cs_n
		inout  wire [15:0] sdram_wire_dq,                    //                          .dq
		output wire [1:0]  sdram_wire_dqm,                   //                          .dqm
		output wire        sdram_wire_ras_n,                 //                          .ras_n
		output wire        sdram_wire_we_n,                  //                          .we_n
		output wire [15:0] second2_export_export,            //            second2_export.export
		output wire [15:0] second_export_export,             //             second_export.export
		output wire [15:0] text_on_export,                   //                   text_on.export
		output wire [15:0] textx_export_export,              //              textx_export.export
		output wire [15:0] texty_export_export,              //              texty_export.export
		output wire [15:0] third2_export_export,             //             third2_export.export
		output wire [15:0] third_export_export               //              third_export.export
	);

	wire         sdram_pll_c0_clk;                                            // sdram_pll:c0 -> [mm_interconnect_0:sdram_pll_c0_clk, rst_controller_001:clk, sdram:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;              // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;               // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                  // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                 // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;             // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire         mm_interconnect_0_text_on_s1_chipselect;                     // mm_interconnect_0:text_on_s1_chipselect -> text_on:chipselect
	wire  [31:0] mm_interconnect_0_text_on_s1_readdata;                       // text_on:readdata -> mm_interconnect_0:text_on_s1_readdata
	wire   [1:0] mm_interconnect_0_text_on_s1_address;                        // mm_interconnect_0:text_on_s1_address -> text_on:address
	wire         mm_interconnect_0_text_on_s1_write;                          // mm_interconnect_0:text_on_s1_write -> text_on:write_n
	wire  [31:0] mm_interconnect_0_text_on_s1_writedata;                      // mm_interconnect_0:text_on_s1_writedata -> text_on:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [1:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_bird_x_s1_chipselect;                      // mm_interconnect_0:bird_x_s1_chipselect -> bird_x:chipselect
	wire  [31:0] mm_interconnect_0_bird_x_s1_readdata;                        // bird_x:readdata -> mm_interconnect_0:bird_x_s1_readdata
	wire   [1:0] mm_interconnect_0_bird_x_s1_address;                         // mm_interconnect_0:bird_x_s1_address -> bird_x:address
	wire         mm_interconnect_0_bird_x_s1_write;                           // mm_interconnect_0:bird_x_s1_write -> bird_x:write_n
	wire  [31:0] mm_interconnect_0_bird_x_s1_writedata;                       // mm_interconnect_0:bird_x_s1_writedata -> bird_x:writedata
	wire         mm_interconnect_0_bird_y_s1_chipselect;                      // mm_interconnect_0:bird_y_s1_chipselect -> bird_y:chipselect
	wire  [31:0] mm_interconnect_0_bird_y_s1_readdata;                        // bird_y:readdata -> mm_interconnect_0:bird_y_s1_readdata
	wire   [1:0] mm_interconnect_0_bird_y_s1_address;                         // mm_interconnect_0:bird_y_s1_address -> bird_y:address
	wire         mm_interconnect_0_bird_y_s1_write;                           // mm_interconnect_0:bird_y_s1_write -> bird_y:write_n
	wire  [31:0] mm_interconnect_0_bird_y_s1_writedata;                       // mm_interconnect_0:bird_y_s1_writedata -> bird_y:writedata
	wire         mm_interconnect_0_pipe1_s1_chipselect;                       // mm_interconnect_0:pipe1_s1_chipselect -> pipe1:chipselect
	wire  [31:0] mm_interconnect_0_pipe1_s1_readdata;                         // pipe1:readdata -> mm_interconnect_0:pipe1_s1_readdata
	wire   [1:0] mm_interconnect_0_pipe1_s1_address;                          // mm_interconnect_0:pipe1_s1_address -> pipe1:address
	wire         mm_interconnect_0_pipe1_s1_write;                            // mm_interconnect_0:pipe1_s1_write -> pipe1:write_n
	wire  [31:0] mm_interconnect_0_pipe1_s1_writedata;                        // mm_interconnect_0:pipe1_s1_writedata -> pipe1:writedata
	wire         mm_interconnect_0_pipe2_s1_chipselect;                       // mm_interconnect_0:pipe2_s1_chipselect -> pipe2:chipselect
	wire  [31:0] mm_interconnect_0_pipe2_s1_readdata;                         // pipe2:readdata -> mm_interconnect_0:pipe2_s1_readdata
	wire   [1:0] mm_interconnect_0_pipe2_s1_address;                          // mm_interconnect_0:pipe2_s1_address -> pipe2:address
	wire         mm_interconnect_0_pipe2_s1_write;                            // mm_interconnect_0:pipe2_s1_write -> pipe2:write_n
	wire  [31:0] mm_interconnect_0_pipe2_s1_writedata;                        // mm_interconnect_0:pipe2_s1_writedata -> pipe2:writedata
	wire         mm_interconnect_0_pipe3_s1_chipselect;                       // mm_interconnect_0:pipe3_s1_chipselect -> pipe3:chipselect
	wire  [31:0] mm_interconnect_0_pipe3_s1_readdata;                         // pipe3:readdata -> mm_interconnect_0:pipe3_s1_readdata
	wire   [1:0] mm_interconnect_0_pipe3_s1_address;                          // mm_interconnect_0:pipe3_s1_address -> pipe3:address
	wire         mm_interconnect_0_pipe3_s1_write;                            // mm_interconnect_0:pipe3_s1_write -> pipe3:write_n
	wire  [31:0] mm_interconnect_0_pipe3_s1_writedata;                        // mm_interconnect_0:pipe3_s1_writedata -> pipe3:writedata
	wire         mm_interconnect_0_pipe_x_s1_chipselect;                      // mm_interconnect_0:pipe_x_s1_chipselect -> pipe_x:chipselect
	wire  [31:0] mm_interconnect_0_pipe_x_s1_readdata;                        // pipe_x:readdata -> mm_interconnect_0:pipe_x_s1_readdata
	wire   [1:0] mm_interconnect_0_pipe_x_s1_address;                         // mm_interconnect_0:pipe_x_s1_address -> pipe_x:address
	wire         mm_interconnect_0_pipe_x_s1_write;                           // mm_interconnect_0:pipe_x_s1_write -> pipe_x:write_n
	wire  [31:0] mm_interconnect_0_pipe_x_s1_writedata;                       // mm_interconnect_0:pipe_x_s1_writedata -> pipe_x:writedata
	wire         mm_interconnect_0_pipe4_s1_chipselect;                       // mm_interconnect_0:pipe4_s1_chipselect -> pipe4:chipselect
	wire  [31:0] mm_interconnect_0_pipe4_s1_readdata;                         // pipe4:readdata -> mm_interconnect_0:pipe4_s1_readdata
	wire   [1:0] mm_interconnect_0_pipe4_s1_address;                          // mm_interconnect_0:pipe4_s1_address -> pipe4:address
	wire         mm_interconnect_0_pipe4_s1_write;                            // mm_interconnect_0:pipe4_s1_write -> pipe4:write_n
	wire  [31:0] mm_interconnect_0_pipe4_s1_writedata;                        // mm_interconnect_0:pipe4_s1_writedata -> pipe4:writedata
	wire         mm_interconnect_0_pipe5_s1_chipselect;                       // mm_interconnect_0:pipe5_s1_chipselect -> pipe5:chipselect
	wire  [31:0] mm_interconnect_0_pipe5_s1_readdata;                         // pipe5:readdata -> mm_interconnect_0:pipe5_s1_readdata
	wire   [1:0] mm_interconnect_0_pipe5_s1_address;                          // mm_interconnect_0:pipe5_s1_address -> pipe5:address
	wire         mm_interconnect_0_pipe5_s1_write;                            // mm_interconnect_0:pipe5_s1_write -> pipe5:write_n
	wire  [31:0] mm_interconnect_0_pipe5_s1_writedata;                        // mm_interconnect_0:pipe5_s1_writedata -> pipe5:writedata
	wire  [31:0] mm_interconnect_0_press_s1_readdata;                         // press:readdata -> mm_interconnect_0:press_s1_readdata
	wire   [1:0] mm_interconnect_0_press_s1_address;                          // mm_interconnect_0:press_s1_address -> press:address
	wire  [31:0] mm_interconnect_0_keycode_s1_readdata;                       // keycode:readdata -> mm_interconnect_0:keycode_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_s1_address;                        // mm_interconnect_0:keycode_s1_address -> keycode:address
	wire         mm_interconnect_0_textx_s1_chipselect;                       // mm_interconnect_0:TextX_s1_chipselect -> TextX:chipselect
	wire  [31:0] mm_interconnect_0_textx_s1_readdata;                         // TextX:readdata -> mm_interconnect_0:TextX_s1_readdata
	wire   [1:0] mm_interconnect_0_textx_s1_address;                          // mm_interconnect_0:TextX_s1_address -> TextX:address
	wire         mm_interconnect_0_textx_s1_write;                            // mm_interconnect_0:TextX_s1_write -> TextX:write_n
	wire  [31:0] mm_interconnect_0_textx_s1_writedata;                        // mm_interconnect_0:TextX_s1_writedata -> TextX:writedata
	wire         mm_interconnect_0_texty_s1_chipselect;                       // mm_interconnect_0:TextY_s1_chipselect -> TextY:chipselect
	wire  [31:0] mm_interconnect_0_texty_s1_readdata;                         // TextY:readdata -> mm_interconnect_0:TextY_s1_readdata
	wire   [1:0] mm_interconnect_0_texty_s1_address;                          // mm_interconnect_0:TextY_s1_address -> TextY:address
	wire         mm_interconnect_0_texty_s1_write;                            // mm_interconnect_0:TextY_s1_write -> TextY:write_n
	wire  [31:0] mm_interconnect_0_texty_s1_writedata;                        // mm_interconnect_0:TextY_s1_writedata -> TextY:writedata
	wire         mm_interconnect_0_first_s1_chipselect;                       // mm_interconnect_0:first_s1_chipselect -> first:chipselect
	wire  [31:0] mm_interconnect_0_first_s1_readdata;                         // first:readdata -> mm_interconnect_0:first_s1_readdata
	wire   [1:0] mm_interconnect_0_first_s1_address;                          // mm_interconnect_0:first_s1_address -> first:address
	wire         mm_interconnect_0_first_s1_write;                            // mm_interconnect_0:first_s1_write -> first:write_n
	wire  [31:0] mm_interconnect_0_first_s1_writedata;                        // mm_interconnect_0:first_s1_writedata -> first:writedata
	wire         mm_interconnect_0_second_s1_chipselect;                      // mm_interconnect_0:second_s1_chipselect -> second:chipselect
	wire  [31:0] mm_interconnect_0_second_s1_readdata;                        // second:readdata -> mm_interconnect_0:second_s1_readdata
	wire   [1:0] mm_interconnect_0_second_s1_address;                         // mm_interconnect_0:second_s1_address -> second:address
	wire         mm_interconnect_0_second_s1_write;                           // mm_interconnect_0:second_s1_write -> second:write_n
	wire  [31:0] mm_interconnect_0_second_s1_writedata;                       // mm_interconnect_0:second_s1_writedata -> second:writedata
	wire         mm_interconnect_0_third_s1_chipselect;                       // mm_interconnect_0:third_s1_chipselect -> third:chipselect
	wire  [31:0] mm_interconnect_0_third_s1_readdata;                         // third:readdata -> mm_interconnect_0:third_s1_readdata
	wire   [1:0] mm_interconnect_0_third_s1_address;                          // mm_interconnect_0:third_s1_address -> third:address
	wire         mm_interconnect_0_third_s1_write;                            // mm_interconnect_0:third_s1_write -> third:write_n
	wire  [31:0] mm_interconnect_0_third_s1_writedata;                        // mm_interconnect_0:third_s1_writedata -> third:writedata
	wire         mm_interconnect_0_scorex_s1_chipselect;                      // mm_interconnect_0:ScoreX_s1_chipselect -> ScoreX:chipselect
	wire  [31:0] mm_interconnect_0_scorex_s1_readdata;                        // ScoreX:readdata -> mm_interconnect_0:ScoreX_s1_readdata
	wire   [1:0] mm_interconnect_0_scorex_s1_address;                         // mm_interconnect_0:ScoreX_s1_address -> ScoreX:address
	wire         mm_interconnect_0_scorex_s1_write;                           // mm_interconnect_0:ScoreX_s1_write -> ScoreX:write_n
	wire  [31:0] mm_interconnect_0_scorex_s1_writedata;                       // mm_interconnect_0:ScoreX_s1_writedata -> ScoreX:writedata
	wire         mm_interconnect_0_scorey_s1_chipselect;                      // mm_interconnect_0:ScoreY_s1_chipselect -> ScoreY:chipselect
	wire  [31:0] mm_interconnect_0_scorey_s1_readdata;                        // ScoreY:readdata -> mm_interconnect_0:ScoreY_s1_readdata
	wire   [1:0] mm_interconnect_0_scorey_s1_address;                         // mm_interconnect_0:ScoreY_s1_address -> ScoreY:address
	wire         mm_interconnect_0_scorey_s1_write;                           // mm_interconnect_0:ScoreY_s1_write -> ScoreY:write_n
	wire  [31:0] mm_interconnect_0_scorey_s1_writedata;                       // mm_interconnect_0:ScoreY_s1_writedata -> ScoreY:writedata
	wire         mm_interconnect_0_scorex2_s1_chipselect;                     // mm_interconnect_0:ScoreX2_s1_chipselect -> ScoreX2:chipselect
	wire  [31:0] mm_interconnect_0_scorex2_s1_readdata;                       // ScoreX2:readdata -> mm_interconnect_0:ScoreX2_s1_readdata
	wire   [1:0] mm_interconnect_0_scorex2_s1_address;                        // mm_interconnect_0:ScoreX2_s1_address -> ScoreX2:address
	wire         mm_interconnect_0_scorex2_s1_write;                          // mm_interconnect_0:ScoreX2_s1_write -> ScoreX2:write_n
	wire  [31:0] mm_interconnect_0_scorex2_s1_writedata;                      // mm_interconnect_0:ScoreX2_s1_writedata -> ScoreX2:writedata
	wire         mm_interconnect_0_scorey2_s1_chipselect;                     // mm_interconnect_0:ScoreY2_s1_chipselect -> ScoreY2:chipselect
	wire  [31:0] mm_interconnect_0_scorey2_s1_readdata;                       // ScoreY2:readdata -> mm_interconnect_0:ScoreY2_s1_readdata
	wire   [1:0] mm_interconnect_0_scorey2_s1_address;                        // mm_interconnect_0:ScoreY2_s1_address -> ScoreY2:address
	wire         mm_interconnect_0_scorey2_s1_write;                          // mm_interconnect_0:ScoreY2_s1_write -> ScoreY2:write_n
	wire  [31:0] mm_interconnect_0_scorey2_s1_writedata;                      // mm_interconnect_0:ScoreY2_s1_writedata -> ScoreY2:writedata
	wire         mm_interconnect_0_bird_y2_s1_chipselect;                     // mm_interconnect_0:bird_y2_s1_chipselect -> bird_y2:chipselect
	wire  [31:0] mm_interconnect_0_bird_y2_s1_readdata;                       // bird_y2:readdata -> mm_interconnect_0:bird_y2_s1_readdata
	wire   [1:0] mm_interconnect_0_bird_y2_s1_address;                        // mm_interconnect_0:bird_y2_s1_address -> bird_y2:address
	wire         mm_interconnect_0_bird_y2_s1_write;                          // mm_interconnect_0:bird_y2_s1_write -> bird_y2:write_n
	wire  [31:0] mm_interconnect_0_bird_y2_s1_writedata;                      // mm_interconnect_0:bird_y2_s1_writedata -> bird_y2:writedata
	wire         mm_interconnect_0_first2_s1_chipselect;                      // mm_interconnect_0:first2_s1_chipselect -> first2:chipselect
	wire  [31:0] mm_interconnect_0_first2_s1_readdata;                        // first2:readdata -> mm_interconnect_0:first2_s1_readdata
	wire   [1:0] mm_interconnect_0_first2_s1_address;                         // mm_interconnect_0:first2_s1_address -> first2:address
	wire         mm_interconnect_0_first2_s1_write;                           // mm_interconnect_0:first2_s1_write -> first2:write_n
	wire  [31:0] mm_interconnect_0_first2_s1_writedata;                       // mm_interconnect_0:first2_s1_writedata -> first2:writedata
	wire         mm_interconnect_0_second2_s1_chipselect;                     // mm_interconnect_0:second2_s1_chipselect -> second2:chipselect
	wire  [31:0] mm_interconnect_0_second2_s1_readdata;                       // second2:readdata -> mm_interconnect_0:second2_s1_readdata
	wire   [1:0] mm_interconnect_0_second2_s1_address;                        // mm_interconnect_0:second2_s1_address -> second2:address
	wire         mm_interconnect_0_second2_s1_write;                          // mm_interconnect_0:second2_s1_write -> second2:write_n
	wire  [31:0] mm_interconnect_0_second2_s1_writedata;                      // mm_interconnect_0:second2_s1_writedata -> second2:writedata
	wire         mm_interconnect_0_third2_s1_chipselect;                      // mm_interconnect_0:third2_s1_chipselect -> third2:chipselect
	wire  [31:0] mm_interconnect_0_third2_s1_readdata;                        // third2:readdata -> mm_interconnect_0:third2_s1_readdata
	wire   [1:0] mm_interconnect_0_third2_s1_address;                         // mm_interconnect_0:third2_s1_address -> third2:address
	wire         mm_interconnect_0_third2_s1_write;                           // mm_interconnect_0:third2_s1_write -> third2:write_n
	wire  [31:0] mm_interconnect_0_third2_s1_writedata;                       // mm_interconnect_0:third2_s1_writedata -> third2:writedata
	wire         mm_interconnect_0_level_s1_chipselect;                       // mm_interconnect_0:level_s1_chipselect -> level:chipselect
	wire  [31:0] mm_interconnect_0_level_s1_readdata;                         // level:readdata -> mm_interconnect_0:level_s1_readdata
	wire   [1:0] mm_interconnect_0_level_s1_address;                          // mm_interconnect_0:level_s1_address -> level:address
	wire         mm_interconnect_0_level_s1_write;                            // mm_interconnect_0:level_s1_write -> level:write_n
	wire  [31:0] mm_interconnect_0_level_s1_writedata;                        // mm_interconnect_0:level_s1_writedata -> level:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [ScoreX2:reset_n, ScoreX:reset_n, ScoreY2:reset_n, ScoreY:reset_n, TextX:reset_n, TextY:reset_n, bird_x:reset_n, bird_y2:reset_n, bird_y:reset_n, first2:reset_n, first:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, keycode:reset_n, level:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, pipe1:reset_n, pipe2:reset_n, pipe3:reset_n, pipe4:reset_n, pipe5:reset_n, pipe_x:reset_n, press:reset_n, rst_translator:in_reset, sdram_pll:reset, second2:reset_n, second:reset_n, sysid_qsys_0:reset_n, text_on:reset_n, third2:reset_n, third:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	flappy_bird_control_ScoreX scorex (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_scorex_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_scorex_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_scorex_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_scorex_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_scorex_s1_readdata),   //                    .readdata
		.out_port   (scorex_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX scorex2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_scorex2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_scorex2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_scorex2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_scorex2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_scorex2_s1_readdata),   //                    .readdata
		.out_port   (scorex2_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX scorey (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_scorey_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_scorey_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_scorey_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_scorey_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_scorey_s1_readdata),   //                    .readdata
		.out_port   (scorey_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX scorey2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_scorey2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_scorey2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_scorey2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_scorey2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_scorey2_s1_readdata),   //                    .readdata
		.out_port   (scorey2_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX textx (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_textx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_textx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_textx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_textx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_textx_s1_readdata),   //                    .readdata
		.out_port   (textx_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX texty (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_texty_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_texty_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_texty_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_texty_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_texty_s1_readdata),   //                    .readdata
		.out_port   (texty_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX bird_x (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_bird_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bird_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bird_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bird_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bird_x_s1_readdata),   //                    .readdata
		.out_port   (bird_x_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX bird_y (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_bird_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bird_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bird_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bird_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bird_y_s1_readdata),   //                    .readdata
		.out_port   (bird_y_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX bird_y2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_bird_y2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bird_y2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bird_y2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bird_y2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bird_y2_s1_readdata),   //                    .readdata
		.out_port   (bird_y2_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX first (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_first_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_first_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_first_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_first_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_first_s1_readdata),   //                    .readdata
		.out_port   (first_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX first2 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_first2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_first2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_first2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_first2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_first2_s1_readdata),   //                    .readdata
		.out_port   (first2_export_export)                    // external_connection.export
	);

	flappy_bird_control_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	flappy_bird_control_keycode keycode (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_keycode_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_keycode_s1_readdata), //                    .readdata
		.in_port  (keycode_export_export)                  // external_connection.export
	);

	flappy_bird_control_ScoreX level (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_level_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_level_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_level_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_level_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_level_s1_readdata),   //                    .readdata
		.out_port   (level_external_connection_export)       // external_connection.export
	);

	flappy_bird_control_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	flappy_bird_control_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	flappy_bird_control_ScoreX pipe1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pipe1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pipe1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pipe1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pipe1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pipe1_s1_readdata),   //                    .readdata
		.out_port   (pipe1_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX pipe2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pipe2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pipe2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pipe2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pipe2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pipe2_s1_readdata),   //                    .readdata
		.out_port   (pipe2_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX pipe3 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pipe3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pipe3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pipe3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pipe3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pipe3_s1_readdata),   //                    .readdata
		.out_port   (pipe3_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX pipe4 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pipe4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pipe4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pipe4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pipe4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pipe4_s1_readdata),   //                    .readdata
		.out_port   (pipe4_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX pipe5 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pipe5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pipe5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pipe5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pipe5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pipe5_s1_readdata),   //                    .readdata
		.out_port   (pipe5_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX pipe_x (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pipe_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pipe_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pipe_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pipe_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pipe_x_s1_readdata),   //                    .readdata
		.out_port   (pipe_x_export_export)                    // external_connection.export
	);

	flappy_bird_control_press press (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_press_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_press_s1_readdata), //                    .readdata
		.in_port  (press_export_export)                  // external_connection.export
	);

	flappy_bird_control_sdram sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	flappy_bird_control_sdram_pll sdram_pll (
		.clk       (clk_clk),                                         //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                  // inclk_interface_reset.reset
		.read      (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0        (sdram_pll_c0_clk),                                //                    c0.clk
		.c1        (sdram_clk_clk),                                   //                    c1.clk
		.areset    (),                                                //        areset_conduit.export
		.locked    (),                                                //        locked_conduit.export
		.phasedone ()                                                 //     phasedone_conduit.export
	);

	flappy_bird_control_ScoreX second (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_second_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_second_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_second_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_second_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_second_s1_readdata),   //                    .readdata
		.out_port   (second_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX second2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_second2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_second2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_second2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_second2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_second2_s1_readdata),   //                    .readdata
		.out_port   (second2_export_export)                    // external_connection.export
	);

	flappy_bird_control_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	flappy_bird_control_ScoreX text_on (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_text_on_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_text_on_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_text_on_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_text_on_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_text_on_s1_readdata),   //                    .readdata
		.out_port   (text_on_export)                           // external_connection.export
	);

	flappy_bird_control_ScoreX third (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_third_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_third_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_third_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_third_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_third_s1_readdata),   //                    .readdata
		.out_port   (third_export_export)                    // external_connection.export
	);

	flappy_bird_control_ScoreX third2 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_third2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_third2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_third2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_third2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_third2_s1_readdata),   //                    .readdata
		.out_port   (third2_export_export)                    // external_connection.export
	);

	flappy_bird_control_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.sdram_pll_c0_clk                               (sdram_pll_c0_clk),                                            //                             sdram_pll_c0.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                          //        sdram_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.bird_x_s1_address                              (mm_interconnect_0_bird_x_s1_address),                         //                                bird_x_s1.address
		.bird_x_s1_write                                (mm_interconnect_0_bird_x_s1_write),                           //                                         .write
		.bird_x_s1_readdata                             (mm_interconnect_0_bird_x_s1_readdata),                        //                                         .readdata
		.bird_x_s1_writedata                            (mm_interconnect_0_bird_x_s1_writedata),                       //                                         .writedata
		.bird_x_s1_chipselect                           (mm_interconnect_0_bird_x_s1_chipselect),                      //                                         .chipselect
		.bird_y_s1_address                              (mm_interconnect_0_bird_y_s1_address),                         //                                bird_y_s1.address
		.bird_y_s1_write                                (mm_interconnect_0_bird_y_s1_write),                           //                                         .write
		.bird_y_s1_readdata                             (mm_interconnect_0_bird_y_s1_readdata),                        //                                         .readdata
		.bird_y_s1_writedata                            (mm_interconnect_0_bird_y_s1_writedata),                       //                                         .writedata
		.bird_y_s1_chipselect                           (mm_interconnect_0_bird_y_s1_chipselect),                      //                                         .chipselect
		.bird_y2_s1_address                             (mm_interconnect_0_bird_y2_s1_address),                        //                               bird_y2_s1.address
		.bird_y2_s1_write                               (mm_interconnect_0_bird_y2_s1_write),                          //                                         .write
		.bird_y2_s1_readdata                            (mm_interconnect_0_bird_y2_s1_readdata),                       //                                         .readdata
		.bird_y2_s1_writedata                           (mm_interconnect_0_bird_y2_s1_writedata),                      //                                         .writedata
		.bird_y2_s1_chipselect                          (mm_interconnect_0_bird_y2_s1_chipselect),                     //                                         .chipselect
		.first_s1_address                               (mm_interconnect_0_first_s1_address),                          //                                 first_s1.address
		.first_s1_write                                 (mm_interconnect_0_first_s1_write),                            //                                         .write
		.first_s1_readdata                              (mm_interconnect_0_first_s1_readdata),                         //                                         .readdata
		.first_s1_writedata                             (mm_interconnect_0_first_s1_writedata),                        //                                         .writedata
		.first_s1_chipselect                            (mm_interconnect_0_first_s1_chipselect),                       //                                         .chipselect
		.first2_s1_address                              (mm_interconnect_0_first2_s1_address),                         //                                first2_s1.address
		.first2_s1_write                                (mm_interconnect_0_first2_s1_write),                           //                                         .write
		.first2_s1_readdata                             (mm_interconnect_0_first2_s1_readdata),                        //                                         .readdata
		.first2_s1_writedata                            (mm_interconnect_0_first2_s1_writedata),                       //                                         .writedata
		.first2_s1_chipselect                           (mm_interconnect_0_first2_s1_chipselect),                      //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.keycode_s1_address                             (mm_interconnect_0_keycode_s1_address),                        //                               keycode_s1.address
		.keycode_s1_readdata                            (mm_interconnect_0_keycode_s1_readdata),                       //                                         .readdata
		.level_s1_address                               (mm_interconnect_0_level_s1_address),                          //                                 level_s1.address
		.level_s1_write                                 (mm_interconnect_0_level_s1_write),                            //                                         .write
		.level_s1_readdata                              (mm_interconnect_0_level_s1_readdata),                         //                                         .readdata
		.level_s1_writedata                             (mm_interconnect_0_level_s1_writedata),                        //                                         .writedata
		.level_s1_chipselect                            (mm_interconnect_0_level_s1_chipselect),                       //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.pipe1_s1_address                               (mm_interconnect_0_pipe1_s1_address),                          //                                 pipe1_s1.address
		.pipe1_s1_write                                 (mm_interconnect_0_pipe1_s1_write),                            //                                         .write
		.pipe1_s1_readdata                              (mm_interconnect_0_pipe1_s1_readdata),                         //                                         .readdata
		.pipe1_s1_writedata                             (mm_interconnect_0_pipe1_s1_writedata),                        //                                         .writedata
		.pipe1_s1_chipselect                            (mm_interconnect_0_pipe1_s1_chipselect),                       //                                         .chipselect
		.pipe2_s1_address                               (mm_interconnect_0_pipe2_s1_address),                          //                                 pipe2_s1.address
		.pipe2_s1_write                                 (mm_interconnect_0_pipe2_s1_write),                            //                                         .write
		.pipe2_s1_readdata                              (mm_interconnect_0_pipe2_s1_readdata),                         //                                         .readdata
		.pipe2_s1_writedata                             (mm_interconnect_0_pipe2_s1_writedata),                        //                                         .writedata
		.pipe2_s1_chipselect                            (mm_interconnect_0_pipe2_s1_chipselect),                       //                                         .chipselect
		.pipe3_s1_address                               (mm_interconnect_0_pipe3_s1_address),                          //                                 pipe3_s1.address
		.pipe3_s1_write                                 (mm_interconnect_0_pipe3_s1_write),                            //                                         .write
		.pipe3_s1_readdata                              (mm_interconnect_0_pipe3_s1_readdata),                         //                                         .readdata
		.pipe3_s1_writedata                             (mm_interconnect_0_pipe3_s1_writedata),                        //                                         .writedata
		.pipe3_s1_chipselect                            (mm_interconnect_0_pipe3_s1_chipselect),                       //                                         .chipselect
		.pipe4_s1_address                               (mm_interconnect_0_pipe4_s1_address),                          //                                 pipe4_s1.address
		.pipe4_s1_write                                 (mm_interconnect_0_pipe4_s1_write),                            //                                         .write
		.pipe4_s1_readdata                              (mm_interconnect_0_pipe4_s1_readdata),                         //                                         .readdata
		.pipe4_s1_writedata                             (mm_interconnect_0_pipe4_s1_writedata),                        //                                         .writedata
		.pipe4_s1_chipselect                            (mm_interconnect_0_pipe4_s1_chipselect),                       //                                         .chipselect
		.pipe5_s1_address                               (mm_interconnect_0_pipe5_s1_address),                          //                                 pipe5_s1.address
		.pipe5_s1_write                                 (mm_interconnect_0_pipe5_s1_write),                            //                                         .write
		.pipe5_s1_readdata                              (mm_interconnect_0_pipe5_s1_readdata),                         //                                         .readdata
		.pipe5_s1_writedata                             (mm_interconnect_0_pipe5_s1_writedata),                        //                                         .writedata
		.pipe5_s1_chipselect                            (mm_interconnect_0_pipe5_s1_chipselect),                       //                                         .chipselect
		.pipe_x_s1_address                              (mm_interconnect_0_pipe_x_s1_address),                         //                                pipe_x_s1.address
		.pipe_x_s1_write                                (mm_interconnect_0_pipe_x_s1_write),                           //                                         .write
		.pipe_x_s1_readdata                             (mm_interconnect_0_pipe_x_s1_readdata),                        //                                         .readdata
		.pipe_x_s1_writedata                            (mm_interconnect_0_pipe_x_s1_writedata),                       //                                         .writedata
		.pipe_x_s1_chipselect                           (mm_interconnect_0_pipe_x_s1_chipselect),                      //                                         .chipselect
		.press_s1_address                               (mm_interconnect_0_press_s1_address),                          //                                 press_s1.address
		.press_s1_readdata                              (mm_interconnect_0_press_s1_readdata),                         //                                         .readdata
		.ScoreX_s1_address                              (mm_interconnect_0_scorex_s1_address),                         //                                ScoreX_s1.address
		.ScoreX_s1_write                                (mm_interconnect_0_scorex_s1_write),                           //                                         .write
		.ScoreX_s1_readdata                             (mm_interconnect_0_scorex_s1_readdata),                        //                                         .readdata
		.ScoreX_s1_writedata                            (mm_interconnect_0_scorex_s1_writedata),                       //                                         .writedata
		.ScoreX_s1_chipselect                           (mm_interconnect_0_scorex_s1_chipselect),                      //                                         .chipselect
		.ScoreX2_s1_address                             (mm_interconnect_0_scorex2_s1_address),                        //                               ScoreX2_s1.address
		.ScoreX2_s1_write                               (mm_interconnect_0_scorex2_s1_write),                          //                                         .write
		.ScoreX2_s1_readdata                            (mm_interconnect_0_scorex2_s1_readdata),                       //                                         .readdata
		.ScoreX2_s1_writedata                           (mm_interconnect_0_scorex2_s1_writedata),                      //                                         .writedata
		.ScoreX2_s1_chipselect                          (mm_interconnect_0_scorex2_s1_chipselect),                     //                                         .chipselect
		.ScoreY_s1_address                              (mm_interconnect_0_scorey_s1_address),                         //                                ScoreY_s1.address
		.ScoreY_s1_write                                (mm_interconnect_0_scorey_s1_write),                           //                                         .write
		.ScoreY_s1_readdata                             (mm_interconnect_0_scorey_s1_readdata),                        //                                         .readdata
		.ScoreY_s1_writedata                            (mm_interconnect_0_scorey_s1_writedata),                       //                                         .writedata
		.ScoreY_s1_chipselect                           (mm_interconnect_0_scorey_s1_chipselect),                      //                                         .chipselect
		.ScoreY2_s1_address                             (mm_interconnect_0_scorey2_s1_address),                        //                               ScoreY2_s1.address
		.ScoreY2_s1_write                               (mm_interconnect_0_scorey2_s1_write),                          //                                         .write
		.ScoreY2_s1_readdata                            (mm_interconnect_0_scorey2_s1_readdata),                       //                                         .readdata
		.ScoreY2_s1_writedata                           (mm_interconnect_0_scorey2_s1_writedata),                      //                                         .writedata
		.ScoreY2_s1_chipselect                          (mm_interconnect_0_scorey2_s1_chipselect),                     //                                         .chipselect
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                          //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                            //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                             //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                         //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                        //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                       //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                      //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                       //                                         .chipselect
		.sdram_pll_pll_slave_address                    (mm_interconnect_0_sdram_pll_pll_slave_address),               //                      sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                      (mm_interconnect_0_sdram_pll_pll_slave_write),                 //                                         .write
		.sdram_pll_pll_slave_read                       (mm_interconnect_0_sdram_pll_pll_slave_read),                  //                                         .read
		.sdram_pll_pll_slave_readdata                   (mm_interconnect_0_sdram_pll_pll_slave_readdata),              //                                         .readdata
		.sdram_pll_pll_slave_writedata                  (mm_interconnect_0_sdram_pll_pll_slave_writedata),             //                                         .writedata
		.second_s1_address                              (mm_interconnect_0_second_s1_address),                         //                                second_s1.address
		.second_s1_write                                (mm_interconnect_0_second_s1_write),                           //                                         .write
		.second_s1_readdata                             (mm_interconnect_0_second_s1_readdata),                        //                                         .readdata
		.second_s1_writedata                            (mm_interconnect_0_second_s1_writedata),                       //                                         .writedata
		.second_s1_chipselect                           (mm_interconnect_0_second_s1_chipselect),                      //                                         .chipselect
		.second2_s1_address                             (mm_interconnect_0_second2_s1_address),                        //                               second2_s1.address
		.second2_s1_write                               (mm_interconnect_0_second2_s1_write),                          //                                         .write
		.second2_s1_readdata                            (mm_interconnect_0_second2_s1_readdata),                       //                                         .readdata
		.second2_s1_writedata                           (mm_interconnect_0_second2_s1_writedata),                      //                                         .writedata
		.second2_s1_chipselect                          (mm_interconnect_0_second2_s1_chipselect),                     //                                         .chipselect
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                         .readdata
		.text_on_s1_address                             (mm_interconnect_0_text_on_s1_address),                        //                               text_on_s1.address
		.text_on_s1_write                               (mm_interconnect_0_text_on_s1_write),                          //                                         .write
		.text_on_s1_readdata                            (mm_interconnect_0_text_on_s1_readdata),                       //                                         .readdata
		.text_on_s1_writedata                           (mm_interconnect_0_text_on_s1_writedata),                      //                                         .writedata
		.text_on_s1_chipselect                          (mm_interconnect_0_text_on_s1_chipselect),                     //                                         .chipselect
		.TextX_s1_address                               (mm_interconnect_0_textx_s1_address),                          //                                 TextX_s1.address
		.TextX_s1_write                                 (mm_interconnect_0_textx_s1_write),                            //                                         .write
		.TextX_s1_readdata                              (mm_interconnect_0_textx_s1_readdata),                         //                                         .readdata
		.TextX_s1_writedata                             (mm_interconnect_0_textx_s1_writedata),                        //                                         .writedata
		.TextX_s1_chipselect                            (mm_interconnect_0_textx_s1_chipselect),                       //                                         .chipselect
		.TextY_s1_address                               (mm_interconnect_0_texty_s1_address),                          //                                 TextY_s1.address
		.TextY_s1_write                                 (mm_interconnect_0_texty_s1_write),                            //                                         .write
		.TextY_s1_readdata                              (mm_interconnect_0_texty_s1_readdata),                         //                                         .readdata
		.TextY_s1_writedata                             (mm_interconnect_0_texty_s1_writedata),                        //                                         .writedata
		.TextY_s1_chipselect                            (mm_interconnect_0_texty_s1_chipselect),                       //                                         .chipselect
		.third_s1_address                               (mm_interconnect_0_third_s1_address),                          //                                 third_s1.address
		.third_s1_write                                 (mm_interconnect_0_third_s1_write),                            //                                         .write
		.third_s1_readdata                              (mm_interconnect_0_third_s1_readdata),                         //                                         .readdata
		.third_s1_writedata                             (mm_interconnect_0_third_s1_writedata),                        //                                         .writedata
		.third_s1_chipselect                            (mm_interconnect_0_third_s1_chipselect),                       //                                         .chipselect
		.third2_s1_address                              (mm_interconnect_0_third2_s1_address),                         //                                third2_s1.address
		.third2_s1_write                                (mm_interconnect_0_third2_s1_write),                           //                                         .write
		.third2_s1_readdata                             (mm_interconnect_0_third2_s1_readdata),                        //                                         .readdata
		.third2_s1_writedata                            (mm_interconnect_0_third2_s1_writedata),                       //                                         .writedata
		.third2_s1_chipselect                           (mm_interconnect_0_third2_s1_chipselect)                       //                                         .chipselect
	);

	flappy_bird_control_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (sdram_pll_c0_clk),                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
